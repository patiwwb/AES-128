--Fichier: InvSbox.vhd
--Auteur: Patryk CHLANDA
--Projet: AES 128 en VHDL
-------
--Copyright 2021, Patryk Chlanda


--imports
library ieee;
use ieee.std_logic_1164.all;
library LIB_AES;
use LIB_AES.state_definition_package.all;

--entity
entity InvSbox is
	port(data_i : in bit8;
	     data_o : out bit8);
end entity;

--architecture
architecture InvSbox_arch of InvSbox is
begin
	--codage de la InvSbox à la main, on peut aussi faire un tableau 
    data_o <= x"63" when data_i = x"00" else
    x"7c" when data_i = x"01" else
    x"77" when data_i = x"02" else
    x"7b" when data_i = x"03" else
    x"f2" when data_i = x"04" else
    x"6b" when data_i = x"05" else
    x"6f" when data_i = x"06" else
    x"c5" when data_i = x"07" else
    x"30" when data_i = x"08" else
    x"01" when data_i = x"09" else
    x"67" when data_i = x"0A" else
    x"2b" when data_i = x"0B" else
    x"fe" when data_i = x"0C" else
    x"d7" when data_i = x"0D" else
    x"ab" when data_i = x"0E" else
    x"76" when data_i = x"0F" else
    x"ca" when data_i = x"10" else
    x"82" when data_i = x"11" else
    x"c9" when data_i = x"12" else
    x"7d" when data_i = x"13" else
    x"fa" when data_i = x"14" else
    x"59" when data_i = x"15" else
    x"47" when data_i = x"16" else
    x"f0" when data_i = x"17" else
    x"ad" when data_i = x"18" else
    x"d4" when data_i = x"19" else
    x"a2" when data_i = x"1A" else
    x"af" when data_i = x"1B" else
    x"9c" when data_i = x"1C" else
    x"a4" when data_i = x"1D" else
    x"72" when data_i = x"1E" else
    x"c0" when data_i = x"1F" else
    x"b7" when data_i = x"20" else
    x"fd" when data_i = x"21" else
    x"93" when data_i = x"22" else
    x"26" when data_i = x"23" else
    x"36" when data_i = x"24" else
    x"3f" when data_i = x"25" else
    x"f7" when data_i = x"26" else
    x"cc" when data_i = x"27" else
    x"34" when data_i = x"28" else
    x"a5" when data_i = x"29" else
    x"e5" when data_i = x"2A" else
    x"f1" when data_i = x"2B" else
    x"71" when data_i = x"2C" else
    x"d8" when data_i = x"2D" else
    x"31" when data_i = x"2E" else
    x"15" when data_i = x"2F" else
    x"04" when data_i = x"30" else
    x"c7" when data_i = x"31" else
    x"23" when data_i = x"32" else
    x"c3" when data_i = x"33" else
    x"18" when data_i = x"34" else
    x"96" when data_i = x"35" else
    x"05" when data_i = x"36" else
    x"9a" when data_i = x"37" else
    x"07" when data_i = x"38" else
    x"12" when data_i = x"39" else
    x"80" when data_i = x"3A" else
    x"e2" when data_i = x"3B" else
    x"eb" when data_i = x"3C" else
    x"27" when data_i = x"3D" else
    x"b2" when data_i = x"3E" else
    x"75" when data_i = x"3F" else
    x"09" when data_i = x"40" else
    x"83" when data_i = x"41" else
    x"2c" when data_i = x"42" else
    x"1a" when data_i = x"43" else
    x"1b" when data_i = x"44" else
    x"6e" when data_i = x"45" else
    x"5a" when data_i = x"46" else
    x"a0" when data_i = x"47" else
    x"52" when data_i = x"48" else
    x"3b" when data_i = x"49" else
    x"d6" when data_i = x"4A" else
    x"b3" when data_i = x"4B" else
    x"29" when data_i = x"4C" else
    x"e3" when data_i = x"4D" else
    x"2f" when data_i = x"4E" else
    x"84" when data_i = x"4F" else
    x"53" when data_i = x"50" else
    x"d1" when data_i = x"51" else
    x"00" when data_i = x"52" else
    x"ed" when data_i = x"53" else
    x"20" when data_i = x"54" else
    x"fc" when data_i = x"55" else
    x"b1" when data_i = x"56" else
    x"5b" when data_i = x"57" else
    x"6a" when data_i = x"58" else
    x"cb" when data_i = x"59" else
    x"be" when data_i = x"5A" else
    x"39" when data_i = x"5B" else
    x"4a" when data_i = x"5C" else
    x"4c" when data_i = x"5D" else
    x"58" when data_i = x"5E" else
    x"cf" when data_i = x"5F" else
    x"d0" when data_i = x"60" else
    x"ef" when data_i = x"61" else
    x"aa" when data_i = x"62" else
    x"fb" when data_i = x"63" else
    x"43" when data_i = x"64" else
    x"4d" when data_i = x"65" else
    x"33" when data_i = x"66" else
    x"85" when data_i = x"67" else
    x"45" when data_i = x"68" else
    x"f9" when data_i = x"69" else
    x"02" when data_i = x"6A" else
    x"7f" when data_i = x"6B" else
    x"50" when data_i = x"6C" else
    x"3c" when data_i = x"6D" else
    x"9f" when data_i = x"6E" else
    x"a8" when data_i = x"6F" else
    x"51" when data_i = x"70" else
    x"a3" when data_i = x"71" else
    x"40" when data_i = x"72" else
    x"8f" when data_i = x"73" else
    x"92" when data_i = x"74" else
    x"9d" when data_i = x"75" else
    x"38" when data_i = x"76" else
    x"f5" when data_i = x"77" else
    x"bc" when data_i = x"78" else
    x"b6" when data_i = x"79" else
    x"da" when data_i = x"7A" else
    x"21" when data_i = x"7B" else
    x"10" when data_i = x"7C" else
    x"ff" when data_i = x"7D" else
    x"f3" when data_i = x"7E" else
    x"d2" when data_i = x"7F" else
    x"cd" when data_i = x"80" else
    x"0c" when data_i = x"81" else
    x"13" when data_i = x"82" else
    x"ec" when data_i = x"83" else
    x"5f" when data_i = x"84" else
    x"97" when data_i = x"85" else
    x"44" when data_i = x"86" else
    x"17" when data_i = x"87" else
    x"c4" when data_i = x"88" else
    x"a7" when data_i = x"89" else
    x"7e" when data_i = x"8A" else
    x"3d" when data_i = x"8B" else
    x"64" when data_i = x"8C" else
    x"5d" when data_i = x"8D" else
    x"19" when data_i = x"8E" else
    x"73" when data_i = x"8F" else
    x"60" when data_i = x"90" else
    x"81" when data_i = x"91" else
    x"4f" when data_i = x"92" else
    x"dc" when data_i = x"93" else
    x"22" when data_i = x"94" else
    x"2a" when data_i = x"95" else
    x"90" when data_i = x"96" else
    x"88" when data_i = x"97" else
    x"46" when data_i = x"98" else
    x"ee" when data_i = x"99" else
    x"b8" when data_i = x"9A" else
    x"14" when data_i = x"9B" else
    x"de" when data_i = x"9C" else
    x"5e" when data_i = x"9D" else
    x"0b" when data_i = x"9E" else
    x"db" when data_i = x"9F" else
    x"e0" when data_i = x"A0" else
    x"32" when data_i = x"A1" else
    x"3a" when data_i = x"A2" else
    x"0a" when data_i = x"A3" else
    x"49" when data_i = x"A4" else
    x"06" when data_i = x"A5" else
    x"24" when data_i = x"A6" else
    x"5c" when data_i = x"A7" else
    x"c2" when data_i = x"A8" else
    x"d3" when data_i = x"A9" else
    x"ac" when data_i = x"AA" else
    x"62" when data_i = x"AB" else
    x"91" when data_i = x"AC" else
    x"95" when data_i = x"AD" else
    x"e4" when data_i = x"AE" else
    x"79" when data_i = x"AF" else
    x"e7" when data_i = x"B0" else
    x"c8" when data_i = x"B1" else
    x"37" when data_i = x"B2" else
    x"6d" when data_i = x"B3" else
    x"8d" when data_i = x"B4" else
    x"d5" when data_i = x"B5" else
    x"4e" when data_i = x"B6" else
    x"a9" when data_i = x"B7" else
    x"6c" when data_i = x"B8" else
    x"56" when data_i = x"B9" else
    x"f4" when data_i = x"BA" else
    x"ea" when data_i = x"BB" else
    x"65" when data_i = x"BC" else
    x"7a" when data_i = x"BD" else
    x"ae" when data_i = x"BE" else
    x"08" when data_i = x"BF" else
    x"ba" when data_i = x"C0" else
    x"78" when data_i = x"C1" else
    x"25" when data_i = x"C2" else
    x"2e" when data_i = x"C3" else
    x"1c" when data_i = x"C4" else
    x"a6" when data_i = x"C5" else
    x"b4" when data_i = x"C6" else
    x"c6" when data_i = x"C7" else
    x"e8" when data_i = x"C8" else
    x"dd" when data_i = x"C9" else
    x"74" when data_i = x"CA" else
    x"1f" when data_i = x"CB" else
    x"4b" when data_i = x"CC" else
    x"bd" when data_i = x"CD" else
    x"8b" when data_i = x"CE" else
    x"8a" when data_i = x"CF" else
    x"70" when data_i = x"D0" else
    x"3e" when data_i = x"D1" else
    x"b5" when data_i = x"D2" else
    x"66" when data_i = x"D3" else
    x"48" when data_i = x"D4" else
    x"03" when data_i = x"D5" else
    x"f6" when data_i = x"D6" else
    x"0e" when data_i = x"D7" else
    x"61" when data_i = x"D8" else
    x"35" when data_i = x"D9" else
    x"57" when data_i = x"DA" else
    x"b9" when data_i = x"DB" else
    x"86" when data_i = x"DC" else
    x"c1" when data_i = x"DD" else
    x"1d" when data_i = x"DE" else
    x"9e" when data_i = x"DF" else
    x"e1" when data_i = x"E0" else
    x"f8" when data_i = x"E1" else
    x"98" when data_i = x"E2" else
    x"11" when data_i = x"E3" else
    x"69" when data_i = x"E4" else
    x"d9" when data_i = x"E5" else
    x"8e" when data_i = x"E6" else
    x"94" when data_i = x"E7" else
    x"9b" when data_i = x"E8" else
    x"1e" when data_i = x"E9" else
    x"87" when data_i = x"EA" else
    x"e9" when data_i = x"EB" else
    x"ce" when data_i = x"EC" else
    x"55" when data_i = x"ED" else
    x"28" when data_i = x"EE" else
    x"df" when data_i = x"EF" else
    x"8c" when data_i = x"F0" else
    x"a1" when data_i = x"F1" else
    x"89" when data_i = x"F2" else
    x"0d" when data_i = x"F3" else
    x"bf" when data_i = x"F4" else
    x"e6" when data_i = x"F5" else
    x"42" when data_i = x"F6" else
    x"68" when data_i = x"F7" else
    x"41" when data_i = x"F8" else
    x"99" when data_i = x"F9" else
    x"2d" when data_i = x"FA" else
    x"0f" when data_i = x"FB" else
    x"b0" when data_i = x"FC" else
    x"54" when data_i = x"FD" else
    x"bb" when data_i = x"FE" else
    x"16" when data_i = x"FF";
	
	
end architecture;
